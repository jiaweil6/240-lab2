`default_nettype none

// ===================
// Submodule Testbench
// ===================

// CompareBlock Testbench

// Subtracter Testbench

// CoinPick Testbench

// UpdateInventory Testbench




// ===================
// Top-level Testbench
// ===================

